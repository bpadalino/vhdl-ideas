package btree is

end package ;
